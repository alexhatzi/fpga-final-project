


module block_module
(
   input wire clk, reset, display_on,
   input wire [9:0] x, y, x_a, y_a,     // current pixel location on screen, without and with arena offset subtracted
   input wire [1:0] cd,                 // bomberman current direction
   input wire [9:0] x_b, y_b,           // bomberman coordinates
   input wire [9:0] waddr,              // write address (a) into block map RAM
   input wire we,                       // write enable to block map RAM
   input wire exp_on,
   output wire [11:0] rgb_out,          // output block rgb
   output wire block_on,                // asserted when x/y within block location on screen
   output wire bm_blocked               // asserted when bomberman is blocked by a block at current location and direction
);

localparam X_WALL_L = 48;                       // end of left wall x coordinate
localparam X_WALL_R = 576;                      // begin of right wall x coordinate
localparam Y_WALL_U = 32;                       // bottom of top wall y coordinate
localparam Y_WALL_D = 448;                      // top of bottom wall y coordinate

localparam BM_HB_OFFSET_9 = 8;                  // offset from top of sprite down to top of 16x16 hit box              
localparam BM_WIDTH       = 16;                 // sprite width
localparam BM_HEIGHT      = 24;                 // sprite height

localparam UP_LEFT_X   = 48;                    // constraints of Bomberman sprite location (upper left corner) within arena.
localparam UP_LEFT_Y   = 32;
localparam LOW_RIGHT_X = 576 - BM_WIDTH;
localparam LOW_RIGHT_Y = 448 - BM_HB_OFFSET_9;    

localparam CD_U = 2'b00;                        // current direction register vals
localparam CD_R = 2'b01;
localparam CD_D = 2'b10;
localparam CD_L = 2'b11;       

// IO for block map dual port RAM
wire data_in = 1'b0; // data input (d)
reg [9:0] raddr;     // read address (dpra)          // write enable (we)
wire data_out;       // data output (dpo)


wire [11:0] dest_out, blk_out ;
reg [3:0] block_dest_state  ;
reg [11:0] dest_animation_addr ; 
reg [26:0] dest_timer ; 
localparam DETS_MAX =  25'd25000000; 

localparam WAIT      = 3'b000 ,
           START     = 3'b001 ,
           FINISH    = 3'b010 ,
           STG1      = 3'b011 ,
           STG2      = 3'b100 , 
           STG3      = 3'b101 , 
           STG4      = 3'b110 , 
           STG5      = 3'b111 ;
             


// signals used to index into block_map RAM to determine if bomberman will collide with a box 
// if moving in a specific direction at the current location. format: <coordinate>_b_hit_<left, right, bottom, top>
wire [9:0] x_b_hit_l, x_b_hit_r, y_b_hit_b, y_b_hit_t;    
wire [9:0] y_b_hit_lr, x_b_hit_bt;

assign x_b_hit_l  = x_b - 1 - X_WALL_L;                   // x coordinate of left  edge of hitbox
assign x_b_hit_r  = x_b + BM_WIDTH - X_WALL_L;            // x coordinate of right edge of hitbox
assign y_b_hit_lr = y_b + BM_HB_OFFSET_9 + 8 - Y_WALL_U;  // y coordinate of middle of hit box

assign y_b_hit_b  = y_b + BM_HEIGHT - Y_WALL_U;           // y coordiante of bottom of hitbox if sprite were going to move down (y + 1)
assign y_b_hit_t  = y_b + BM_HB_OFFSET_9 - 1 - Y_WALL_U;  // y coordinate of top of hitbox if sprite were going to move up (y - 1)
assign x_b_hit_bt = x_b + 7 - X_WALL_L;                   // x coordinate of middle of hitbox

// read address into block_map RAM
// first address condition reads into RAM for current ABM coordinate of VGA pixel on screen to display blocks
// next four address conditions index into RAM to check block_map if a block is in bomberman's path to assert bm_blocked output           
always @(posedge clk)
   begin
   if(display_on & x > X_WALL_L & x < X_WALL_R & y > Y_WALL_U & y < Y_WALL_D+16)
      raddr = x_a[9:4] + y_a[9:4]*33;
   else if(!display_on)
      begin
      if(cd == CD_L)
         raddr = x_b_hit_l[9:4]  + y_b_hit_lr[9:4]*33;
      else if(cd == CD_R)
         raddr = x_b_hit_r[9:4]  + y_b_hit_lr[9:4]*33;
      else if(cd == CD_U)
         raddr = x_b_hit_bt[9:4] +  y_b_hit_t[9:4]*33;
      else 
         raddr = x_b_hit_bt[9:4] +  y_b_hit_b[9:4]*33;
      end
   else 
      raddr = 896; // don't care index in RAM
   end


   always @ ( posedge clk ) begin
      case (block_dest_state)
      WAIT : begin
               if (block_on & exp_on ) 
               block_dest_state <= START ; 
              end
      START : begin
               dest_animation_addr <= (x_a[3:0]) + {(y_a[3:0]), 4'd0} ; 
                  if (dest_timer == DETS_MAX ) begin
                     dest_timer <= 0 ; 
                     block_dest_state <= STG1 ; 
                  end else dest_timer <= dest_timer + 1 ; 
              end      
      STG1 : begin
               dest_animation_addr <= (x_a[3:0]) + {(y_a[3:0]), 4'd0} + 256  ; 
                  if (dest_timer == DETS_MAX ) begin
                     dest_timer <= 0 ; 
                     block_dest_state <= STG2 ; 
                  end else dest_timer <= dest_timer + 1 ; 
              end      
      STG2 : begin
               dest_animation_addr <= (x_a[3:0]) + {(y_a[3:0]), 4'd0} + 512 ; 
                  if (dest_timer == DETS_MAX ) begin
                     dest_timer <= 0 ; 
                     block_dest_state <= STG3 ; 
                  end else dest_timer <= dest_timer + 1 ; 
              end      
      STG3 : begin
               dest_animation_addr <= (x_a[3:0]) + {(y_a[3:0]), 4'd0} +  768 ; 
                  if (dest_timer == DETS_MAX ) begin
                     dest_timer <= 0 ; 
                     block_dest_state <= STG4 ; 
                  end else dest_timer <= dest_timer + 1 ; 
              end      
      STG4 : begin
               dest_animation_addr <= (x_a[3:0]) + {(y_a[3:0]), 4'd0} + 1024 ; 
                  if (dest_timer == DETS_MAX ) begin
                     dest_timer <= 0 ; 
                     block_dest_state <= STG5 ; 
                  end else dest_timer <= dest_timer + 1 ; 
              end      
      STG5 : begin
               dest_animation_addr <= (x_a[3:0]) + {(y_a[3:0]), 4'd0} + 1280 ; 
                  if (dest_timer == DETS_MAX ) begin
                     dest_timer <= 0 ; 
                     block_dest_state <= FINISH ; 
                  end else dest_timer <= dest_timer + 1 ; 
              end      
      FINISH : begin
                 block_dest_state <= WAIT  ;
              end      

      endcase
   end


// instantiate block sprite ROM
// index into ROM uses x/y pixel arena coordinates lower 4 bits, as each block is 16x16
block_dm block_unit(.a((x_a[3:0]) + {(y_a[3:0]), 4'd0}), .spo(blk_out));
block_dest_rom block_dest_unit (.a(dest_animation_addr), .spo(dest_out)) ; 

// instantiate block_map distributed dual port RAM
block_map block_map_unit(.a(waddr), .d(data_in), .dpra(raddr), .clk(clk), .we(we), .spo(), .dpo(data_out));
   
// register to hold state of bomberman being blocked in current direction by a block
reg blocked_reg; 
wire blocked_next;

always @(posedge clk, posedge reset)
   if(reset)
      blocked_reg <= 0;
   else 
      blocked_reg <= blocked_next;
      
assign rgb_out   = (exp_on & block_on) ? dest_out : blk_out ; 

// check output of block_map when !display_on and raddr is looking for a block in bomberman's path
assign blocked_next = (!display_on & data_out == 1) ? 1 : 
                      (!display_on & data_out == 0) ? 0 : blocked_reg;

// assert when bomberman is blocked by a block
assign bm_blocked = blocked_reg;

// assert when display is on and output from block_map is 1, indicating x/y is in a block
assign block_on = display_on & data_out; 

endmodule
